-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Fri Dec 05 11:33:13 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY timerNEANDER IS 
	PORT
	(
		reset :  IN  STD_LOGIC;
		clock :  IN  STD_LOGIC;
		goto_t0 :  IN  STD_LOGIC;
		t :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END timerNEANDER;

ARCHITECTURE bdf_type OF timerNEANDER IS 

COMPONENT mux4p1
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 Sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 S : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	and0t1 :  STD_LOGIC;
SIGNAL	and0t2 :  STD_LOGIC;
SIGNAL	and0t3 :  STD_LOGIC;
SIGNAL	clock_real :  STD_LOGIC;
SIGNAL	D :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	not_w :  STD_LOGIC;
SIGNAL	or1 :  STD_LOGIC;
SIGNAL	or2 :  STD_LOGIC;
SIGNAL	or3 :  STD_LOGIC;
SIGNAL	Sel :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	t_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	w :  STD_LOGIC;
SIGNAL	x :  STD_LOGIC;
SIGNAL	y :  STD_LOGIC;
SIGNAL	z :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;


BEGIN 



and0t2 <= and0t1 AND z;



and0t1 <= x AND y;


PROCESS(clock_real,reset)
BEGIN
IF (reset = '0') THEN
	x <= '0';
ELSIF (RISING_EDGE(clock_real)) THEN
	x <= SYNTHESIZED_WIRE_0;
END IF;
END PROCESS;


PROCESS(clock_real,reset)
BEGIN
IF (reset = '0') THEN
	y <= '0';
ELSIF (RISING_EDGE(clock_real)) THEN
	y <= SYNTHESIZED_WIRE_1;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_18 <= NOT(x);



SYNTHESIZED_WIRE_16 <= NOT(z);



t_ALTERA_SYNTHESIZED(2) <= SYNTHESIZED_WIRE_2 AND SYNTHESIZED_WIRE_3 AND y AND not_w;


t_ALTERA_SYNTHESIZED(3) <= x AND SYNTHESIZED_WIRE_4 AND y AND not_w;


SYNTHESIZED_WIRE_31 <= NOT(y);



SYNTHESIZED_WIRE_30 <= NOT(z);



SYNTHESIZED_WIRE_2 <= NOT(x);



t_ALTERA_SYNTHESIZED(4) <= SYNTHESIZED_WIRE_5 AND z AND SYNTHESIZED_WIRE_6 AND not_w;


SYNTHESIZED_WIRE_3 <= NOT(z);



t_ALTERA_SYNTHESIZED(5) <= x AND z AND SYNTHESIZED_WIRE_7 AND not_w;



SYNTHESIZED_WIRE_4 <= NOT(z);



SYNTHESIZED_WIRE_5 <= NOT(x);



SYNTHESIZED_WIRE_6 <= NOT(y);



t_ALTERA_SYNTHESIZED(6) <= SYNTHESIZED_WIRE_8 AND z AND y AND not_w;


t_ALTERA_SYNTHESIZED(7) <= x AND z AND y AND not_w;


SYNTHESIZED_WIRE_7 <= NOT(y);



SYNTHESIZED_WIRE_8 <= NOT(x);



SYNTHESIZED_WIRE_20 <= NOT(y);




Sel(1) <= NOT(goto_t0);



PROCESS(clock_real,reset)
BEGIN
IF (reset = '0') THEN
	z <= '0';
ELSIF (RISING_EDGE(clock_real)) THEN
	z <= SYNTHESIZED_WIRE_9;
END IF;
END PROCESS;


PROCESS(clock_real,reset)
BEGIN
IF (reset = '0') THEN
	w <= '0';
ELSIF (RISING_EDGE(clock_real)) THEN
	w <= SYNTHESIZED_WIRE_10;
END IF;
END PROCESS;


b2v_inst31 : mux4p1
PORT MAP(A => D(2),
		 B => z,
		 C => SYNTHESIZED_WIRE_11,
		 D => SYNTHESIZED_WIRE_12,
		 Sel => Sel,
		 S => SYNTHESIZED_WIRE_9);


b2v_inst32 : mux4p1
PORT MAP(A => D(3),
		 B => w,
		 C => SYNTHESIZED_WIRE_13,
		 D => SYNTHESIZED_WIRE_14,
		 Sel => Sel,
		 S => SYNTHESIZED_WIRE_10);


SYNTHESIZED_WIRE_19 <= NOT(z);



SYNTHESIZED_WIRE_22 <= NOT(y);



SYNTHESIZED_WIRE_21 <= NOT(z);



SYNTHESIZED_WIRE_23 <= NOT(x);



SYNTHESIZED_WIRE_24 <= NOT(z);



SYNTHESIZED_WIRE_25 <= NOT(z);



SYNTHESIZED_WIRE_26 <= NOT(x);



t_ALTERA_SYNTHESIZED(0) <= SYNTHESIZED_WIRE_15 AND SYNTHESIZED_WIRE_16 AND SYNTHESIZED_WIRE_17 AND not_w;


SYNTHESIZED_WIRE_27 <= NOT(y);



SYNTHESIZED_WIRE_28 <= NOT(y);



SYNTHESIZED_WIRE_29 <= NOT(x);



t_ALTERA_SYNTHESIZED(8) <= SYNTHESIZED_WIRE_18 AND SYNTHESIZED_WIRE_19 AND SYNTHESIZED_WIRE_20 AND w;


t_ALTERA_SYNTHESIZED(9) <= x AND SYNTHESIZED_WIRE_21 AND SYNTHESIZED_WIRE_22 AND w;


t_ALTERA_SYNTHESIZED(10) <= SYNTHESIZED_WIRE_23 AND SYNTHESIZED_WIRE_24 AND y AND w;


t_ALTERA_SYNTHESIZED(11) <= x AND SYNTHESIZED_WIRE_25 AND y AND w;


t_ALTERA_SYNTHESIZED(12) <= SYNTHESIZED_WIRE_26 AND z AND SYNTHESIZED_WIRE_27 AND w;


t_ALTERA_SYNTHESIZED(13) <= x AND z AND SYNTHESIZED_WIRE_28 AND w;


t_ALTERA_SYNTHESIZED(14) <= SYNTHESIZED_WIRE_29 AND z AND y AND w;


t_ALTERA_SYNTHESIZED(1) <= x AND SYNTHESIZED_WIRE_30 AND SYNTHESIZED_WIRE_31 AND not_w;


t_ALTERA_SYNTHESIZED(15) <= x AND z AND y AND w;


not_w <= NOT(w);



SYNTHESIZED_WIRE_15 <= NOT(x);



SYNTHESIZED_WIRE_38 <= NOT(SYNTHESIZED_WIRE_39);



SYNTHESIZED_WIRE_12 <= NOT(SYNTHESIZED_WIRE_33);



SYNTHESIZED_WIRE_14 <= NOT(SYNTHESIZED_WIRE_34);



SYNTHESIZED_WIRE_17 <= NOT(y);



b2v_inst8 : mux4p1
PORT MAP(A => D(0),
		 B => x,
		 C => SYNTHESIZED_WIRE_40,
		 D => SYNTHESIZED_WIRE_40,
		 Sel => Sel,
		 S => SYNTHESIZED_WIRE_0);


b2v_inst9 : mux4p1
PORT MAP(A => D(1),
		 B => y,
		 C => SYNTHESIZED_WIRE_39,
		 D => SYNTHESIZED_WIRE_38,
		 Sel => Sel,
		 S => SYNTHESIZED_WIRE_1);


SYNTHESIZED_WIRE_40 <= NOT(x);



or1 <= y OR x;


or2 <= z OR or1;



SYNTHESIZED_WIRE_11 <= z XOR and0t1;


SYNTHESIZED_WIRE_13 <= w XOR and0t2;


SYNTHESIZED_WIRE_39 <= y XOR x;


SYNTHESIZED_WIRE_33 <= z XOR or1;


SYNTHESIZED_WIRE_34 <= w XOR or2;

t <= t_ALTERA_SYNTHESIZED;
clock_real <= clock;

Sel(0) <= '0';
END bdf_type;