-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Wed Dec 17 03:22:45 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY decoderNEANDER IS 
	PORT
	(
		clk :  IN  STD_LOGIC;
		Nflag :  IN  STD_LOGIC;
		Zflag :  IN  STD_LOGIC;
		A :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		CargaPC :  OUT  STD_LOGIC;
		CargaREM :  OUT  STD_LOGIC;
		IncrementaPC :  OUT  STD_LOGIC;
		CargaRI :  OUT  STD_LOGIC;
		sel_literalmente_so_sel :  OUT  STD_LOGIC;
		CargaRDM :  OUT  STD_LOGIC;
		Read :  OUT  STD_LOGIC;
		Write :  OUT  STD_LOGIC;
		CargaAC :  OUT  STD_LOGIC;
		CargaNZ :  OUT  STD_LOGIC;
		halted :  OUT  STD_LOGIC;
		ULAencoder :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END decoderNEANDER;

ARCHITECTURE bdf_type OF decoderNEANDER IS 

COMPONENT timerneander
	PORT(goto_t0 : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 t : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	ADD :  STD_LOGIC;
SIGNAL	ANDx :  STD_LOGIC;
SIGNAL	goto_t0 :  STD_LOGIC;
SIGNAL	HLT :  STD_LOGIC;
SIGNAL	JMP :  STD_LOGIC;
SIGNAL	JN :  STD_LOGIC;
SIGNAL	JUMP_CONFIRMADO :  STD_LOGIC;
SIGNAL	JZ :  STD_LOGIC;
SIGNAL	LDA :  STD_LOGIC;
SIGNAL	NEG :  STD_LOGIC;
SIGNAL	NOP :  STD_LOGIC;
SIGNAL	NOTx :  STD_LOGIC;
SIGNAL	ORx :  STD_LOGIC;
SIGNAL	STA :  STD_LOGIC;
SIGNAL	SUB :  STD_LOGIC;
SIGNAL	t :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	ULA_COM_OPERANDO :  STD_LOGIC;
SIGNAL	ULA_SEM_OPERANDO :  STD_LOGIC;
SIGNAL	ULAencoder_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	XORx :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;


BEGIN 
CargaAC <= SYNTHESIZED_WIRE_67;
CargaNZ <= SYNTHESIZED_WIRE_67;
SYNTHESIZED_WIRE_13 <= '1';



sel_literalmente_so_sel <= t(7) AND SYNTHESIZED_WIRE_0;


STA <= SYNTHESIZED_WIRE_68 AND SYNTHESIZED_WIRE_69 AND SYNTHESIZED_WIRE_70 AND A(0);


HLT <= A(3) AND A(2) AND A(1) AND A(0);


ULA_SEM_OPERANDO <= NOTx OR NEG;


XORx <= SYNTHESIZED_WIRE_68 AND A(2) AND A(1) AND A(0);


NEG <= A(3) AND A(2) AND SYNTHESIZED_WIRE_70 AND SYNTHESIZED_WIRE_71;


SUB <= A(3) AND A(2) AND SYNTHESIZED_WIRE_70 AND A(0);


SYNTHESIZED_WIRE_22 <= JN AND Nflag;


SYNTHESIZED_WIRE_9 <= SUB OR ANDx OR ADD;


SYNTHESIZED_WIRE_8 <= XORx OR LDA OR ORx;


ULA_COM_OPERANDO <= SYNTHESIZED_WIRE_8 OR SYNTHESIZED_WIRE_9;



LDA <= SYNTHESIZED_WIRE_68 AND SYNTHESIZED_WIRE_69 AND A(1) AND SYNTHESIZED_WIRE_71;


b2v_inst20 : timerneander
PORT MAP(goto_t0 => goto_t0,
		 reset => SYNTHESIZED_WIRE_13,
		 clock => clk,
		 t => t);


SYNTHESIZED_WIRE_71 <= NOT(A(0));



SYNTHESIZED_WIRE_70 <= NOT(A(1));



SYNTHESIZED_WIRE_69 <= NOT(A(2));



SYNTHESIZED_WIRE_68 <= NOT(A(3));



SYNTHESIZED_WIRE_17 <= NOT(HLT);



SYNTHESIZED_WIRE_23 <= JZ AND Zflag;


goto_t0 <= SYNTHESIZED_WIRE_14 OR SYNTHESIZED_WIRE_15 OR HLT OR SYNTHESIZED_WIRE_16;


SYNTHESIZED_WIRE_34 <= SYNTHESIZED_WIRE_17 AND t(1);


ADD <= SYNTHESIZED_WIRE_68 AND SYNTHESIZED_WIRE_69 AND A(1) AND A(0);


CargaREM <= SYNTHESIZED_WIRE_20 AND SYNTHESIZED_WIRE_21;


SYNTHESIZED_WIRE_20 <= NOT(HLT);



JUMP_CONFIRMADO <= SYNTHESIZED_WIRE_22 OR JMP OR SYNTHESIZED_WIRE_23;


CargaPC <= JUMP_CONFIRMADO AND t(7);


CargaRI <= SYNTHESIZED_WIRE_24 AND t(3);


SYNTHESIZED_WIRE_24 <= NOT(HLT);



ORx <= SYNTHESIZED_WIRE_68 AND A(2) AND SYNTHESIZED_WIRE_70 AND SYNTHESIZED_WIRE_71;


SYNTHESIZED_WIRE_21 <= SYNTHESIZED_WIRE_28 OR SYNTHESIZED_WIRE_29 OR t(0);


SYNTHESIZED_WIRE_28 <= t(4) AND SYNTHESIZED_WIRE_30;


SYNTHESIZED_WIRE_30 <= STA OR JUMP_CONFIRMADO OR ULA_COM_OPERANDO;


SYNTHESIZED_WIRE_29 <= t(7) AND SYNTHESIZED_WIRE_31;


SYNTHESIZED_WIRE_31 <= STA OR ULA_COM_OPERANDO;


IncrementaPC <= SYNTHESIZED_WIRE_32 OR SYNTHESIZED_WIRE_33 OR SYNTHESIZED_WIRE_34;


ANDx <= SYNTHESIZED_WIRE_68 AND A(2) AND SYNTHESIZED_WIRE_70 AND A(0);


SYNTHESIZED_WIRE_32 <= SYNTHESIZED_WIRE_37 AND t(4);


SYNTHESIZED_WIRE_37 <= STA OR ULA_COM_OPERANDO;


SYNTHESIZED_WIRE_33 <= t(3) AND SYNTHESIZED_WIRE_38;


SYNTHESIZED_WIRE_42 <= SYNTHESIZED_WIRE_39 AND JN;


SYNTHESIZED_WIRE_41 <= SYNTHESIZED_WIRE_40 AND JZ;


SYNTHESIZED_WIRE_38 <= SYNTHESIZED_WIRE_41 OR SYNTHESIZED_WIRE_42;


SYNTHESIZED_WIRE_39 <= NOT(Nflag);



SYNTHESIZED_WIRE_40 <= NOT(Zflag);



SYNTHESIZED_WIRE_0 <= STA OR ULA_COM_OPERANDO;


NOTx <= SYNTHESIZED_WIRE_68 AND A(2) AND A(1) AND SYNTHESIZED_WIRE_71;


CargaRDM <= t(9) AND STA;


Read <= SYNTHESIZED_WIRE_45 OR SYNTHESIZED_WIRE_46 OR t(2);


SYNTHESIZED_WIRE_45 <= t(6) AND SYNTHESIZED_WIRE_47;


SYNTHESIZED_WIRE_47 <= STA OR JUMP_CONFIRMADO OR ULA_COM_OPERANDO;


SYNTHESIZED_WIRE_46 <= t(9) AND ULA_COM_OPERANDO;


Write <= t(10) AND STA;


ULAencoder_ALTERA_SYNTHESIZED(0) <= NEG AND t(4);


ULAencoder_ALTERA_SYNTHESIZED(1) <= SUB AND t(10);


ULAencoder_ALTERA_SYNTHESIZED(2) <= LDA AND t(10);


JMP <= A(3) AND SYNTHESIZED_WIRE_69 AND SYNTHESIZED_WIRE_70 AND SYNTHESIZED_WIRE_71;


ULAencoder_ALTERA_SYNTHESIZED(3) <= ADD AND t(10);


ULAencoder_ALTERA_SYNTHESIZED(4) <= ORx AND t(10);


ULAencoder_ALTERA_SYNTHESIZED(5) <= ANDx AND t(10);


ULAencoder_ALTERA_SYNTHESIZED(6) <= NOTx AND t(4);


ULAencoder_ALTERA_SYNTHESIZED(7) <= XORx AND t(10);


SYNTHESIZED_WIRE_51 <= ULA_COM_OPERANDO AND t(10);


SYNTHESIZED_WIRE_67 <= SYNTHESIZED_WIRE_51 OR SYNTHESIZED_WIRE_52;


SYNTHESIZED_WIRE_52 <= ULA_SEM_OPERANDO AND t(4);


SYNTHESIZED_WIRE_14 <= t(10) AND SYNTHESIZED_WIRE_53;


JN <= A(3) AND SYNTHESIZED_WIRE_69 AND SYNTHESIZED_WIRE_70 AND A(0);


SYNTHESIZED_WIRE_53 <= STA OR ULA_COM_OPERANDO;


SYNTHESIZED_WIRE_16 <= t(4) AND SYNTHESIZED_WIRE_56;


SYNTHESIZED_WIRE_56 <= NOP OR SYNTHESIZED_WIRE_57 OR SYNTHESIZED_WIRE_58 OR ULA_SEM_OPERANDO;


SYNTHESIZED_WIRE_57 <= JZ AND SYNTHESIZED_WIRE_59;


SYNTHESIZED_WIRE_58 <= JN AND SYNTHESIZED_WIRE_60;


SYNTHESIZED_WIRE_59 <= NOT(Zflag);



SYNTHESIZED_WIRE_60 <= NOT(Nflag);



SYNTHESIZED_WIRE_15 <= t(7) AND JUMP_CONFIRMADO;


JZ <= A(3) AND SYNTHESIZED_WIRE_69 AND A(1) AND SYNTHESIZED_WIRE_71;


NOP <= SYNTHESIZED_WIRE_68 AND SYNTHESIZED_WIRE_69 AND SYNTHESIZED_WIRE_70 AND SYNTHESIZED_WIRE_71;

halted <= HLT;
ULAencoder <= ULAencoder_ALTERA_SYNTHESIZED;

END bdf_type;