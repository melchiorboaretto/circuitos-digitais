-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Tue Nov 25 22:49:49 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY program_counter IS 
	PORT
	(
		reset :  IN  STD_LOGIC;
		clock :  IN  STD_LOGIC;
		D :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		Sel :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		S :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END program_counter;

ARCHITECTURE bdf_type OF program_counter IS 

COMPONENT mux4p1
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 Sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 S : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	and0t1 :  STD_LOGIC;
SIGNAL	and0t2 :  STD_LOGIC;
SIGNAL	and0t3 :  STD_LOGIC;
SIGNAL	and0t4 :  STD_LOGIC;
SIGNAL	and0t5 :  STD_LOGIC;
SIGNAL	and0t6 :  STD_LOGIC;
SIGNAL	clock_real :  STD_LOGIC;
SIGNAL	or1 :  STD_LOGIC;
SIGNAL	or2 :  STD_LOGIC;
SIGNAL	or3 :  STD_LOGIC;
SIGNAL	or4 :  STD_LOGIC;
SIGNAL	or5 :  STD_LOGIC;
SIGNAL	or6 :  STD_LOGIC;
SIGNAL	S_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;


BEGIN 



and0t2 <= and0t1 AND S_ALTERA_SYNTHESIZED(2);


and0t3 <= and0t2 AND S_ALTERA_SYNTHESIZED(3);


and0t4 <= and0t3 AND S_ALTERA_SYNTHESIZED(4);


and0t5 <= and0t4 AND S_ALTERA_SYNTHESIZED(5);


and0t6 <= and0t5 AND S_ALTERA_SYNTHESIZED(6);


and0t1 <= S_ALTERA_SYNTHESIZED(0) AND S_ALTERA_SYNTHESIZED(1);


PROCESS(clock_real,reset)
BEGIN
IF (reset = '0') THEN
	S_ALTERA_SYNTHESIZED(0) <= '0';
ELSIF (RISING_EDGE(clock_real)) THEN
	S_ALTERA_SYNTHESIZED(0) <= SYNTHESIZED_WIRE_0;
END IF;
END PROCESS;


PROCESS(clock_real,reset)
BEGIN
IF (reset = '0') THEN
	S_ALTERA_SYNTHESIZED(1) <= '0';
ELSIF (RISING_EDGE(clock_real)) THEN
	S_ALTERA_SYNTHESIZED(1) <= SYNTHESIZED_WIRE_1;
END IF;
END PROCESS;


b2v_inst10 : mux4p1
PORT MAP(A => D(2),
		 B => S_ALTERA_SYNTHESIZED(2),
		 C => SYNTHESIZED_WIRE_2,
		 D => SYNTHESIZED_WIRE_3,
		 Sel => Sel,
		 S => SYNTHESIZED_WIRE_14);


b2v_inst11 : mux4p1
PORT MAP(A => D(3),
		 B => S_ALTERA_SYNTHESIZED(3),
		 C => SYNTHESIZED_WIRE_4,
		 D => SYNTHESIZED_WIRE_5,
		 Sel => Sel,
		 S => SYNTHESIZED_WIRE_15);


b2v_inst12 : mux4p1
PORT MAP(A => D(4),
		 B => S_ALTERA_SYNTHESIZED(4),
		 C => SYNTHESIZED_WIRE_6,
		 D => SYNTHESIZED_WIRE_7,
		 Sel => Sel,
		 S => SYNTHESIZED_WIRE_16);


b2v_inst13 : mux4p1
PORT MAP(A => D(5),
		 B => S_ALTERA_SYNTHESIZED(5),
		 C => SYNTHESIZED_WIRE_8,
		 D => SYNTHESIZED_WIRE_9,
		 Sel => Sel,
		 S => SYNTHESIZED_WIRE_17);


b2v_inst14 : mux4p1
PORT MAP(A => D(6),
		 B => S_ALTERA_SYNTHESIZED(6),
		 C => SYNTHESIZED_WIRE_10,
		 D => SYNTHESIZED_WIRE_11,
		 Sel => Sel,
		 S => SYNTHESIZED_WIRE_18);


b2v_inst15 : mux4p1
PORT MAP(A => D(7),
		 B => S_ALTERA_SYNTHESIZED(7),
		 C => SYNTHESIZED_WIRE_12,
		 D => SYNTHESIZED_WIRE_13,
		 Sel => Sel,
		 S => SYNTHESIZED_WIRE_26);


PROCESS(clock_real,reset)
BEGIN
IF (reset = '0') THEN
	S_ALTERA_SYNTHESIZED(2) <= '0';
ELSIF (RISING_EDGE(clock_real)) THEN
	S_ALTERA_SYNTHESIZED(2) <= SYNTHESIZED_WIRE_14;
END IF;
END PROCESS;


PROCESS(clock_real,reset)
BEGIN
IF (reset = '0') THEN
	S_ALTERA_SYNTHESIZED(3) <= '0';
ELSIF (RISING_EDGE(clock_real)) THEN
	S_ALTERA_SYNTHESIZED(3) <= SYNTHESIZED_WIRE_15;
END IF;
END PROCESS;


PROCESS(clock_real,reset)
BEGIN
IF (reset = '0') THEN
	S_ALTERA_SYNTHESIZED(4) <= '0';
ELSIF (RISING_EDGE(clock_real)) THEN
	S_ALTERA_SYNTHESIZED(4) <= SYNTHESIZED_WIRE_16;
END IF;
END PROCESS;


PROCESS(clock_real,reset)
BEGIN
IF (reset = '0') THEN
	S_ALTERA_SYNTHESIZED(5) <= '0';
ELSIF (RISING_EDGE(clock_real)) THEN
	S_ALTERA_SYNTHESIZED(5) <= SYNTHESIZED_WIRE_17;
END IF;
END PROCESS;


PROCESS(clock_real,reset)
BEGIN
IF (reset = '0') THEN
	S_ALTERA_SYNTHESIZED(6) <= '0';
ELSIF (RISING_EDGE(clock_real)) THEN
	S_ALTERA_SYNTHESIZED(6) <= SYNTHESIZED_WIRE_18;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_30 <= NOT(SYNTHESIZED_WIRE_31);



SYNTHESIZED_WIRE_3 <= NOT(SYNTHESIZED_WIRE_20);



SYNTHESIZED_WIRE_5 <= NOT(SYNTHESIZED_WIRE_21);



SYNTHESIZED_WIRE_7 <= NOT(SYNTHESIZED_WIRE_22);



SYNTHESIZED_WIRE_9 <= NOT(SYNTHESIZED_WIRE_23);



SYNTHESIZED_WIRE_11 <= NOT(SYNTHESIZED_WIRE_24);



SYNTHESIZED_WIRE_13 <= NOT(SYNTHESIZED_WIRE_25);



PROCESS(clock_real,reset)
BEGIN
IF (reset = '0') THEN
	S_ALTERA_SYNTHESIZED(7) <= '0';
ELSIF (RISING_EDGE(clock_real)) THEN
	S_ALTERA_SYNTHESIZED(7) <= SYNTHESIZED_WIRE_26;
END IF;
END PROCESS;


b2v_inst8 : mux4p1
PORT MAP(A => D(0),
		 B => S_ALTERA_SYNTHESIZED(0),
		 C => SYNTHESIZED_WIRE_32,
		 D => SYNTHESIZED_WIRE_32,
		 Sel => Sel,
		 S => SYNTHESIZED_WIRE_0);


b2v_inst9 : mux4p1
PORT MAP(A => D(1),
		 B => S_ALTERA_SYNTHESIZED(1),
		 C => SYNTHESIZED_WIRE_31,
		 D => SYNTHESIZED_WIRE_30,
		 Sel => Sel,
		 S => SYNTHESIZED_WIRE_1);


SYNTHESIZED_WIRE_32 <= NOT(S_ALTERA_SYNTHESIZED(0));



or1 <= S_ALTERA_SYNTHESIZED(1) OR S_ALTERA_SYNTHESIZED(0);


or2 <= S_ALTERA_SYNTHESIZED(2) OR or1;


or3 <= S_ALTERA_SYNTHESIZED(3) OR or2;


or4 <= S_ALTERA_SYNTHESIZED(4) OR or3;


or5 <= S_ALTERA_SYNTHESIZED(5) OR or4;


or6 <= S_ALTERA_SYNTHESIZED(6) OR or5;


SYNTHESIZED_WIRE_2 <= S_ALTERA_SYNTHESIZED(2) XOR and0t1;


SYNTHESIZED_WIRE_4 <= S_ALTERA_SYNTHESIZED(3) XOR and0t2;


SYNTHESIZED_WIRE_6 <= S_ALTERA_SYNTHESIZED(4) XOR and0t3;


SYNTHESIZED_WIRE_8 <= S_ALTERA_SYNTHESIZED(5) XOR and0t4;


SYNTHESIZED_WIRE_10 <= S_ALTERA_SYNTHESIZED(6) XOR and0t5;


SYNTHESIZED_WIRE_12 <= S_ALTERA_SYNTHESIZED(7) XOR and0t6;


SYNTHESIZED_WIRE_31 <= S_ALTERA_SYNTHESIZED(1) XOR S_ALTERA_SYNTHESIZED(0);


SYNTHESIZED_WIRE_20 <= S_ALTERA_SYNTHESIZED(2) XOR or1;


SYNTHESIZED_WIRE_21 <= S_ALTERA_SYNTHESIZED(3) XOR or2;


SYNTHESIZED_WIRE_22 <= S_ALTERA_SYNTHESIZED(4) XOR or3;


SYNTHESIZED_WIRE_23 <= S_ALTERA_SYNTHESIZED(5) XOR or4;


SYNTHESIZED_WIRE_24 <= S_ALTERA_SYNTHESIZED(6) XOR or5;


SYNTHESIZED_WIRE_25 <= S_ALTERA_SYNTHESIZED(7) XOR or6;

S <= S_ALTERA_SYNTHESIZED;
clock_real <= clock;

END bdf_type;