-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Tue Nov 25 00:37:04 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY ula8bNEANDER IS 
	PORT
	(
		A :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		B :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		opSel :  IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
		N :  OUT  STD_LOGIC;
		Z :  OUT  STD_LOGIC;
		S :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END ula8bNEANDER;

ARCHITECTURE bdf_type OF ula8bNEANDER IS 

COMPONENT mux8b8
	PORT(A : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 C : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 D : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 E : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 F : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 G : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 H : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 Sel : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 S : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT cslaclas8
	PORT(sel : IN STD_LOGIC;
		 A : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 Cout : OUT STD_LOGIC;
		 S : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT signinv8b
	PORT(E : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 S : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT tap8
	PORT(Barramento : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 S0 : OUT STD_LOGIC;
		 S1 : OUT STD_LOGIC;
		 S2 : OUT STD_LOGIC;
		 S3 : OUT STD_LOGIC;
		 S4 : OUT STD_LOGIC;
		 S5 : OUT STD_LOGIC;
		 S6 : OUT STD_LOGIC;
		 S7 : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	N_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	S_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;


BEGIN 



b2v_inst : mux8b8
PORT MAP(A => SYNTHESIZED_WIRE_22,
		 B => SYNTHESIZED_WIRE_1,
		 C => SYNTHESIZED_WIRE_2,
		 D => SYNTHESIZED_WIRE_3,
		 E => SYNTHESIZED_WIRE_4,
		 F => SYNTHESIZED_WIRE_5,
		 G => SYNTHESIZED_WIRE_22,
		 H => B,
		 Sel => opSel,
		 S => S_ALTERA_SYNTHESIZED);


SYNTHESIZED_WIRE_1 <= A AND B;


Z <= SYNTHESIZED_WIRE_7 AND SYNTHESIZED_WIRE_8 AND SYNTHESIZED_WIRE_9 AND SYNTHESIZED_WIRE_10 AND SYNTHESIZED_WIRE_11 AND SYNTHESIZED_WIRE_12 AND SYNTHESIZED_WIRE_13 AND SYNTHESIZED_WIRE_14;


SYNTHESIZED_WIRE_14 <= NOT(SYNTHESIZED_WIRE_15);



SYNTHESIZED_WIRE_9 <= NOT(SYNTHESIZED_WIRE_16);



SYNTHESIZED_WIRE_12 <= NOT(SYNTHESIZED_WIRE_17);



SYNTHESIZED_WIRE_10 <= NOT(SYNTHESIZED_WIRE_18);



SYNTHESIZED_WIRE_11 <= NOT(SYNTHESIZED_WIRE_19);



SYNTHESIZED_WIRE_13 <= NOT(N_ALTERA_SYNTHESIZED);



SYNTHESIZED_WIRE_2 <= B OR A;


SYNTHESIZED_WIRE_3 <= NOT(A);



b2v_inst4 : cslaclas8
PORT MAP(sel => opSel(2),
		 A => A,
		 B => B,
		 S => SYNTHESIZED_WIRE_22);


b2v_inst5 : signinv8b
PORT MAP(E => A,
		 S => SYNTHESIZED_WIRE_5);


SYNTHESIZED_WIRE_4 <= A XOR B;


SYNTHESIZED_WIRE_7 <= NOT(SYNTHESIZED_WIRE_20);



SYNTHESIZED_WIRE_8 <= NOT(SYNTHESIZED_WIRE_21);



b2v_inst9 : tap8
PORT MAP(Barramento => S_ALTERA_SYNTHESIZED,
		 S0 => SYNTHESIZED_WIRE_20,
		 S1 => SYNTHESIZED_WIRE_16,
		 S2 => SYNTHESIZED_WIRE_21,
		 S3 => SYNTHESIZED_WIRE_18,
		 S4 => SYNTHESIZED_WIRE_15,
		 S5 => SYNTHESIZED_WIRE_17,
		 S6 => SYNTHESIZED_WIRE_19,
		 S7 => N_ALTERA_SYNTHESIZED);

N <= N_ALTERA_SYNTHESIZED;
S <= S_ALTERA_SYNTHESIZED;

END bdf_type;