-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Wed Dec 03 17:41:49 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY decoderNEANDER IS 
	PORT
	(
		clk :  IN  STD_LOGIC;
		Nflag :  IN  STD_LOGIC;
		Zflag :  IN  STD_LOGIC;
		A :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		CargaPC :  OUT  STD_LOGIC;
		CargaREM :  OUT  STD_LOGIC;
		IncrementaPC :  OUT  STD_LOGIC;
		CargaRI :  OUT  STD_LOGIC;
		sel_literalmente_so_sel :  OUT  STD_LOGIC;
		CargaRDM :  OUT  STD_LOGIC;
		Read :  OUT  STD_LOGIC;
		Write :  OUT  STD_LOGIC;
		CargaAC :  OUT  STD_LOGIC;
		CargaNZ :  OUT  STD_LOGIC;
		ULAencoder :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END decoderNEANDER;

ARCHITECTURE bdf_type OF decoderNEANDER IS 

COMPONENT timerneander
	PORT(goto_t0 : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 t : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	ADD :  STD_LOGIC;
SIGNAL	ANDx :  STD_LOGIC;
SIGNAL	goto_t0 :  STD_LOGIC;
SIGNAL	HLT :  STD_LOGIC;
SIGNAL	JMP :  STD_LOGIC;
SIGNAL	JN :  STD_LOGIC;
SIGNAL	JUMP_CONFIRMADO :  STD_LOGIC;
SIGNAL	JZ :  STD_LOGIC;
SIGNAL	LDA :  STD_LOGIC;
SIGNAL	NEG :  STD_LOGIC;
SIGNAL	NOP :  STD_LOGIC;
SIGNAL	NOTx :  STD_LOGIC;
SIGNAL	ORx :  STD_LOGIC;
SIGNAL	STA :  STD_LOGIC;
SIGNAL	SUB :  STD_LOGIC;
SIGNAL	t :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	ULA_COM_OPERANDO :  STD_LOGIC;
SIGNAL	ULA_SEM_OPERANDO :  STD_LOGIC;
SIGNAL	ULAencoder_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	XORx :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;


BEGIN 
CargaAC <= SYNTHESIZED_WIRE_62;
CargaNZ <= SYNTHESIZED_WIRE_62;
SYNTHESIZED_WIRE_17 <= '1';



sel_literalmente_so_sel <= t(5) AND SYNTHESIZED_WIRE_0;


STA <= SYNTHESIZED_WIRE_63 AND SYNTHESIZED_WIRE_64 AND SYNTHESIZED_WIRE_65 AND A(0);



ULA_SEM_OPERANDO <= NOTx OR NEG;


XORx <= SYNTHESIZED_WIRE_63 AND A(2) AND A(1) AND A(0);


NEG <= A(3) AND A(2) AND SYNTHESIZED_WIRE_65 AND SYNTHESIZED_WIRE_66;


SUB <= A(3) AND A(2) AND SYNTHESIZED_WIRE_65 AND A(0);


SYNTHESIZED_WIRE_15 <= JN AND Nflag;


SYNTHESIZED_WIRE_9 <= SUB OR ANDx OR ADD;


SYNTHESIZED_WIRE_8 <= XORx OR LDA OR ORx;


ULA_COM_OPERANDO <= SYNTHESIZED_WIRE_8 OR SYNTHESIZED_WIRE_9;



LDA <= SYNTHESIZED_WIRE_63 AND SYNTHESIZED_WIRE_64 AND A(1) AND SYNTHESIZED_WIRE_66;


SYNTHESIZED_WIRE_66 <= NOT(A(0));



SYNTHESIZED_WIRE_65 <= NOT(A(1));



SYNTHESIZED_WIRE_64 <= NOT(A(2));



SYNTHESIZED_WIRE_63 <= NOT(A(3));



SYNTHESIZED_WIRE_16 <= JZ AND Zflag;


ADD <= SYNTHESIZED_WIRE_63 AND SYNTHESIZED_WIRE_64 AND A(1) AND A(0);


JUMP_CONFIRMADO <= SYNTHESIZED_WIRE_15 OR JMP OR SYNTHESIZED_WIRE_16;


CargaPC <= JUMP_CONFIRMADO AND t(5);


b2v_inst39 : timerneander
PORT MAP(goto_t0 => goto_t0,
		 reset => SYNTHESIZED_WIRE_17,
		 clock => clk,
		 t => t);


ORx <= SYNTHESIZED_WIRE_63 AND A(2) AND SYNTHESIZED_WIRE_65 AND SYNTHESIZED_WIRE_66;


CargaREM <= SYNTHESIZED_WIRE_21 OR SYNTHESIZED_WIRE_22 OR t(0);


SYNTHESIZED_WIRE_21 <= t(3) AND SYNTHESIZED_WIRE_23;


SYNTHESIZED_WIRE_23 <= STA OR JUMP_CONFIRMADO OR ULA_COM_OPERANDO;


SYNTHESIZED_WIRE_22 <= t(5) AND SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_24 <= STA OR ULA_COM_OPERANDO;


IncrementaPC <= SYNTHESIZED_WIRE_25 OR SYNTHESIZED_WIRE_26 OR t(1);


ANDx <= SYNTHESIZED_WIRE_63 AND A(2) AND SYNTHESIZED_WIRE_65 AND A(0);


SYNTHESIZED_WIRE_25 <= SYNTHESIZED_WIRE_29 AND t(4);


SYNTHESIZED_WIRE_29 <= STA OR ULA_COM_OPERANDO;


SYNTHESIZED_WIRE_26 <= t(3) AND SYNTHESIZED_WIRE_30;


SYNTHESIZED_WIRE_34 <= SYNTHESIZED_WIRE_31 AND JN;


SYNTHESIZED_WIRE_33 <= SYNTHESIZED_WIRE_32 AND JZ;


SYNTHESIZED_WIRE_30 <= SYNTHESIZED_WIRE_33 OR SYNTHESIZED_WIRE_34;


SYNTHESIZED_WIRE_31 <= NOT(Nflag);



SYNTHESIZED_WIRE_32 <= NOT(Zflag);



SYNTHESIZED_WIRE_0 <= STA OR ULA_COM_OPERANDO;


NOTx <= SYNTHESIZED_WIRE_63 AND A(2) AND A(1) AND SYNTHESIZED_WIRE_66;


CargaRDM <= t(6) AND STA;


Read <= SYNTHESIZED_WIRE_37 OR SYNTHESIZED_WIRE_38 OR t(1);


SYNTHESIZED_WIRE_37 <= t(4) AND SYNTHESIZED_WIRE_39;


SYNTHESIZED_WIRE_39 <= STA OR JUMP_CONFIRMADO OR ULA_COM_OPERANDO;


SYNTHESIZED_WIRE_38 <= t(6) AND ULA_COM_OPERANDO;


Write <= t(7) AND STA;


ULAencoder_ALTERA_SYNTHESIZED(0) <= NEG AND t(3);


ULAencoder_ALTERA_SYNTHESIZED(1) <= SUB AND t(7);


ULAencoder_ALTERA_SYNTHESIZED(2) <= LDA AND t(7);


JMP <= A(3) AND SYNTHESIZED_WIRE_64 AND SYNTHESIZED_WIRE_65 AND SYNTHESIZED_WIRE_66;


ULAencoder_ALTERA_SYNTHESIZED(3) <= ADD AND t(7);


ULAencoder_ALTERA_SYNTHESIZED(4) <= ORx AND t(7);


ULAencoder_ALTERA_SYNTHESIZED(5) <= ANDx AND t(7);


ULAencoder_ALTERA_SYNTHESIZED(6) <= NOTx AND t(3);


ULAencoder_ALTERA_SYNTHESIZED(7) <= XORx AND t(7);


SYNTHESIZED_WIRE_43 <= ULA_COM_OPERANDO AND t(7);


SYNTHESIZED_WIRE_62 <= SYNTHESIZED_WIRE_43 OR SYNTHESIZED_WIRE_44;


SYNTHESIZED_WIRE_44 <= ULA_SEM_OPERANDO AND t(3);


SYNTHESIZED_WIRE_50 <= t(7) AND SYNTHESIZED_WIRE_45;


JN <= A(3) AND SYNTHESIZED_WIRE_64 AND SYNTHESIZED_WIRE_65 AND A(0);


SYNTHESIZED_WIRE_45 <= STA OR ULA_COM_OPERANDO;


goto_t0 <= SYNTHESIZED_WIRE_48 OR SYNTHESIZED_WIRE_49 OR SYNTHESIZED_WIRE_50;


SYNTHESIZED_WIRE_48 <= t(3) AND SYNTHESIZED_WIRE_51;


SYNTHESIZED_WIRE_51 <= NOP OR SYNTHESIZED_WIRE_52 OR SYNTHESIZED_WIRE_53 OR ULA_SEM_OPERANDO;


SYNTHESIZED_WIRE_52 <= JZ AND SYNTHESIZED_WIRE_54;


SYNTHESIZED_WIRE_53 <= JN AND SYNTHESIZED_WIRE_55;


SYNTHESIZED_WIRE_54 <= NOT(Zflag);



SYNTHESIZED_WIRE_55 <= NOT(Nflag);



SYNTHESIZED_WIRE_49 <= t(5) AND JUMP_CONFIRMADO;


JZ <= A(3) AND SYNTHESIZED_WIRE_64 AND A(1) AND SYNTHESIZED_WIRE_66;


NOP <= SYNTHESIZED_WIRE_63 AND SYNTHESIZED_WIRE_64 AND SYNTHESIZED_WIRE_65 AND SYNTHESIZED_WIRE_66;

CargaRI <= t(2);
ULAencoder <= ULAencoder_ALTERA_SYNTHESIZED;

END bdf_type;